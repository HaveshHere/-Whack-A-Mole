module BoardTest(input wire [3:0]sw, output wire [3:0]LEDR);

   assign LEDR = sw;
	
endmodule
